//  Top-level processor module

module processor (
			     );

// Skeleton
		
// Instantiate Program counter register
// PC+4
// Shift left 26
// Control unit after decoding --> forward nets to mux's and alu
// RegFile
// Sign extender
// ALU control
// ALU
// Shift left 32
// Adder
// Memory

// Mux's as we go

// Considerations: Reordering of modules to reduce clock cycles

endmodule